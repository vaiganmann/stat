library verilog;
use verilog.vl_types.all;
entity definitions_main is
end definitions_main;
