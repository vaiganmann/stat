library verilog;
use verilog.vl_types.all;
entity definitions is
end definitions;
