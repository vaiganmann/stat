library verilog;
use verilog.vl_types.all;
entity definitions_bus is
end definitions_bus;
