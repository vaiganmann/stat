library verilog;
use verilog.vl_types.all;
entity definitions_mem is
end definitions_mem;
